---------------------------------------------------------------------------
-- program_counter.vhd - Program Counter Implementation 
-- 
-- Note : The program counter is simply a register that updates its output 
-- on the rising clock edge.
-- 
--
-- Copyright (C) 2006 by Lih Wen Koh (lwkoh@cse.unsw.edu.au)
-- All Rights Reserved. 
--
-- The single-cycle processor core is provided AS IS, with no warranty of 
-- any kind, express or implied. The user of the program accepts full 
-- responsibility for the application of the program and the use of any 
-- results. This work may be downloaded, compiled, executed, copied, and 
-- modified solely for nonprofit, educational, noncommercial research, and 
-- noncommercial scholarship purposes provided that this notice in its 
-- entirety accompanies all copies. Copies of the modified software can be 
-- delivered to persons who use it solely for nonprofit, educational, 
-- noncommercial research, and noncommercial scholarship purposes provided 
-- that this notice in its entirety accompanies all copies.
--
---------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity program_counter is
    port ( reset    : in  std_logic;
           stall    : in std_logic;
           clk      : in  std_logic;
           addr_in  : in  std_logic_vector(3 downto 0);
           addr_out : out std_logic_vector(3 downto 0) );
end program_counter;

architecture behavioral of program_counter is
begin

    update_process: process ( reset, 
                              clk ) is
    begin
        if (falling_edge(clk)) then
            if (stall = '0') then
                addr_out <= addr_in;
            end if; 
        end if;
        
        if (falling_edge(reset)) then
           addr_out <= (others => '0'); 
        end if;

    end process;
end behavioral;
